
`define registers_addr_width 4
`define registers_data_width 32
